-- Katie Pucci
-- COE1502:: CPU
-- Forwarding Control Unit

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY forwarding_unit IS
    -- Define ports
    -- Inputs::
    --
    -- Outputs::
    --
    PORT (

    );

END forwarding_unit;

ARCHITECTURE Behavioral OF forwarding_unit IS

BEGIN

    PROCESS ()
    BEGIN

    END PROCESS;



END Behavioral;
